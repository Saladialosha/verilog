module btgtb();
reg b0,b1,b2,b3;
wire g0,g1,g2,g3;
btg m3(b0,b1,b2,b3,g0,g1,g2,g3);
initial
begin
b3=0; b2=0; b1=0; b0=0;
#2
b3=0; b2=0; b1=0; b0=1;
#2
b3=0; b2=0; b1=1; b0=0;
#2
b3=0; b2=0; b1=1; b0=1;
#2
b3=0; b2=1; b1=0; b0=0;
#2
b3=0; b2=1; b1=0; b0=1;
#2
b3=0; b2=1; b1=1; b0=0;
#2
b3=0; b2=1; b1=1; b0=1;
#2
b3=1; b2=0; b1=0; b0=0;
#2
b3=1; b2=0; b1=0; b0=1;
#2
b3=1; b2=0; b1=1; b0=0;
#2
b3=1; b2=0; b1=1; b0=1;
#2
b3=1; b2=1; b1=0; b0=0;
#2
b3=1; b2=1; b1=0; b0=1;
#2
b3=1; b2=1; b1=1; b0=0;
#2
b3=1; b2=1; b1=1; b0=1;
#5 $stop;
end
endmodule
